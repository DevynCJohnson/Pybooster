[styling]
attribute=attribute
block_comment=block_comment
comment=comment
comment_line_bang=comment_line_bang
identifier=identifier
keyword=keyword
number=number
operator=operator
stdfunction=stdfunction
stdoperator=stdoperator
stdpackage=stdpackage
stdtype=stdtype
string=string
stringeol=stringeol
userword=type

[keywords]
attributes=active ascending base delayed driving driving_value event high image instance_name last_active last_event last_value left leftof length low path_name pos pred quiet range reverse_range right rightof simple_name stable succ transaction val value
docComment=a addindex addtogroup anchor annotatedclasslist arg attention author authors b brief bug c callergraph callgraph category cite class classhierarchy code cond copybrief copydetails copydoc copyright date def defgroup define deprecated details diafile dir docbookonly dontinclude dot dotfile e else elseif em endcode endcond enddocbookonly enddot endhtmlonly endif endinternal endlatexonly endlink endmanonly endmsc endparblock endrtfonly endsecreflist enduml endverbatim endxmlonly enum example exception extends ff[ f] file fn functionindex f{ f} header headerfile headerfilelist hidecallergraph hidecallgraph hideinitializer htmlinclude htmlonly idlexcept if ifnot image implements include includedoc includelineno ingroup inherit interface internal invariant l latexinclude latexonly li license line link mainpage manonly memberof msc mscfile n name namespace nosubgrouping note overload p package page par paragraph param param[in] parblock post postheader pre private privatesection property protected protectedsection protocol public publicsection pure ref refitem related relatedalso relates relatesalso remark remarks result return returns retval rtfonly sa secreflist section see short showinitializer since skip skipline snippet snippetdoc snippetlineno startuml static struct subpage subsection subsubsection tableofcontents test throw throws todo tparam typedef union until var verbatim verbinclude version vhdlflow warning weakgroup xmlonly xrefitem
keywords=access after alias all architecture array assert attribute begin block body buffer bus case component configuration constant disconnect downto else elsif end entity exit file for function generate generic group guarded if impure in inertial inout is label library linkage literal loop map new next null of on open others out package port postponed procedure process pure range record register reject report return select severity shared signal subtype then to transport type unaffected units until use variable wait when while with
operators=abs and mod nand nor not or rem rol ror sla sll sra srl xnor xor
std_functions=endfile falling_edge is_x now read readline resize resolved rising_edge rotate_left rotate_right shift_left shift_right std_match to_01 to_bit to_bitvector to_integer to_signed to_stdlogicvector to_stdulogic to_stdulogicvector to_unsigned to_UX01 to_x01 to_x01z write writeline
std_packages=ieee math_complex math_real numeric_bit numeric_std standard std std_logic_1164 std_logic_arith std_logic_misc std_logic_signed std_logic_textio std_logic_unsigned textio vital_primitives vital_timing work
std_types=bit bit_vector boolean character delay_length file_open_kind file_open_status integer line natural positive real severity_level side signed std_logic std_logic_vector std_ulogic std_ulogic_vector string text time unsigned UX01 UX01Z width X01 X01Z
userwords=

[lexer_properties]
fold.at.Begin=1
fold.at.else=1
fold.at.Parenthese=1
fold.at.When=1
fold.comment=1
fold.compact=0

[settings]
extension=vhd
mime_type=text/x-vhdl
comment_single=--
comment_use_indent=true
context_action_cmd=

[indentation]
type=1
width=4
